��C      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�K �min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G?޸Q���feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Oxygen��Temperature��Humidity�et�b�n_features_in_�K�
n_outputs_�K�classes_�hhK ��h��R�(KK��h �i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���h4C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��h4�C       �t�bK��R�}�(h	K�
node_count�K�nodes�hhK ��h��R�(KK��h �V56�����R�(Kh$N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hVh4K ��hWh4K��hXh4K��hYh �f8�����R�(Kh5NNNJ����J����K t�bK��hZhdK ��h[h4K(��h\hdK0��uK8KKt�b�C�                         ���?�G�z��?<             N@������������������������       �                     ;@������������������������       �        !            �@@�t�b�values�hhK ��h��R�(KKKK��hd�C0      ;@     �@@      ;@                     �@@�t�bub�_sklearn_version��1.1.2�ub.
����      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.2�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG?��G�z�feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Oxygen��Temperature��Humidity�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��h2�f8�����R�(KhGNNNJ����J����K t�b�C              �?�t�bhKh&�scalar���hFC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK�
node_count�K�nodes�h(h+K ��h-��R�(KK��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hwhFK ��hxhFK��hyhFK��hzhWK��h{hWK ��h|hFK(��h}hWK0��uK8KKt�b�C�                        p���?      �?&             N@������������������������       �ȵHPS!�?             :@������������������������       �H�V�e��?             A@�t�b�values�h(h+K ��h-��R�(KKKK��hW�C0      >@      >@      @      7@      ;@      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ��g�?�G�z��?(             N@������������������������       �                     ;@������������������������       �                    �@@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ;@     �@@      ;@                     �@@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?��Q��?$             N@������������������������       �                     5@������������������������       �                    �C@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      5@     �C@      5@                     �C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?*;L]n�?%             N@������������������������       �@4և���?             <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@       @              @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         �Y7�?��S���?)             N@������������������������       �                     @@������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      @@      <@      @@                      <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�0u��A�?'             N@������������������������       �                     7@������������������������       �                    �B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      7@     �B@      7@                     �B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��������?$             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      =@      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?      �?'             N@������������������������       �      �?             @@������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      >@      >@      >@       @              <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?*;L]n�?)             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         �|��?*;L]n�?"             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJQY%hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�G�z��?$             N@������������������������       �                    �@@������������������������       �                     ;@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0     �@@      ;@     �@@                      ;@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��fbhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�0u��A�?'             N@������������������������       �                     7@������������������������       �                    �B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      7@     �B@      7@                     �B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$�phG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ���0u���?&             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      1@     �E@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW:+LhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ���Q��?%             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      5@     �C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF<KdhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?d��0u��?#             N@������������������������       �                     6@������������������������       �                     C@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      6@      C@      6@                      C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJؽ�hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��G�z��?(             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      ;@     �@@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJX��vhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�q�q�?(             N@������������������������       �                     9@������������������������       �                    �A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      9@     �A@      9@                     �A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���EhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?�G�z��?'             N@������������������������       �                     ;@������������������������       �                    �@@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ;@     �@@      ;@                     �@@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:9)bhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�������?&             N@������������������������       �(;L]n�?             >@������������������������       �                     >@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      =@      �?              >@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�BHzhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?�������?%             N@������������������������       �                     =@������������������������       �                     ?@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      =@                      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�}�JhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��������?(             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      =@      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ'J�OhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?*;L]n�?(             N@������������������������       �                     A@������������������������       �                     :@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      A@      :@      A@                      :@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW�ehG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ��g�?��S���?,             N@������������������������       �                     <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      <@      @@      <@                      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���zhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?�G�z��?(             N@������������������������       �                    �@@������������������������       �                     ;@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0     �@@      ;@     �@@                      ;@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJX^khG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?*;L]n�?(             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJQ��dhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?��S���?!             N@������������������������       �                     @@������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      @@      <@      @@                      <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���lhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?�q�q�?&             N@������������������������       �                     9@������������������������       �                    �A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      9@     �A@      9@                     �A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJB	VhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��������?#             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      ?@      =@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJMk/hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��q�q�?'             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C     �A@      9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJH�_VhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?*;L]n�?$             N@������������������������       �                     A@������������������������       �                     :@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      A@      :@      A@                      :@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	NhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?*;L]n�?(             N@������������������������       �                     9@������������������������       ���?^�k�?            �A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      9@              �?      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���%hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ���S���?%             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      @@      <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJs-hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        0I��?�0u��A�?&             N@������������������������       �                     7@������������������������       �                    �B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      7@     �B@      7@                     �B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�E^hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?�q�q�?%             N@������������������������       �                    �A@������������������������       �                     9@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0     �A@      9@     �A@                      9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�&UhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�������?%             N@������������������������       �                     <@������������������������       �      �?             @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      <@              �?      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�uhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�B                          `!�?�G�z��?$             N@������������������������       �P���Q�?             4@                        �$I�?��Q��?             D@������������������������       �                     :@������������������������       �        	             ,@�t�bh�h(h+K ��h-��R�(KKKK��hW�CP      ;@     �@@      �?      3@      :@      ,@      :@                      ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�G5GhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?�������?&             N@������������������������       �                     ?@������������������������       �                     =@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ?@      =@      ?@                      =@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJO�#hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�G�z��?)             N@������������������������       �                    �@@������������������������       �                     ;@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0     �@@      ;@     �@@                      ;@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��^hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?*;L]n�?#             N@������������������������       �                     7@������������������������       ��L���?            �B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      7@              @      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�	�^hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ���S���?)             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      <@      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJR��zhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?*;L]n�?(             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJc`>yhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�B                          ���?��Q��?(             N@                        ����?�+e�X�?"             I@������������������������       �        
             (@������������������������       �                     C@������������������������       �ףp=
�?             $@�t�bh�h(h+K ��h-��R�(KKKK��hW�CP      5@     �C@      (@      C@      (@                      C@      "@      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJا�LhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�G�z��?&             N@������������������������       �h�����?             <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ;@     �@@      ;@      �?              @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�|MhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?�������?#             N@������������������������       �                     ?@������������������������       �                     =@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ?@      =@      ?@                      =@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�#vhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       �d��0u��?&             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      6@      C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ>hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?��S���?%             N@������������������������       �                     <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      <@      @@      <@                      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���GhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?���Q��?'             N@������������������������       �                     8@������������������������       �                     B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      8@      B@      8@                      B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��-hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?*;L]n�?*             N@������������������������       �                    �@@������������������������       � 7���B�?             ;@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      A@      :@     �@@              �?      :@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�;GhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?���Q��?&             N@������������������������       �                     8@������������������������       �                     B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      8@      B@      8@                      B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�a{8hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�q�q�?#             N@������������������������       �                     9@������������������������       �                    �A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      9@     �A@      9@                     �A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ ��#hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �\;�?*;L]n�?%             N@������������������������       �:�&���?            �C@������������������������       ������?             5@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      @      @@      3@       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�?�hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?*;L]n�?'             N@������������������������       �                     8@������������������������       ��X�<ݺ?             B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      8@               @      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	Ͳ$hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�������?$             N@������������������������       �      �?             @@������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ?@      =@      ?@      �?              <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�J�	hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        0I��?�q�q�?$             N@������������������������       �                     9@������������������������       �                    �A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      9@     �A@      9@                     �A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��qhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �m��?�������?(             N@������������������������       �(;L]n�?             >@������������������������       �                     >@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      =@      �?              >@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ �4BhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ��g�?��S���?'             N@������������������������       �                     <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      <@      @@      <@                      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJڗhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�G�z��?)             N@������������������������       � 	��p�?             =@������������������������       �                     ?@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ;@     �@@      ;@       @              ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       �*;L]n�?(             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      :@      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�H'jhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��q�q�?%             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      9@     �A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��=yhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�q�q�?$             N@������������������������       � �Cc}�?             <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      9@     �A@      9@      @              @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��ChG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         �|��?���Q��?)             N@������������������������       �                     8@������������������������       �                     B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      8@      B@      8@                      B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�y�/hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?���Q��?%             N@������������������������       �                     6@������������������������       ��}�+r��?             C@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      8@      B@      6@               @      B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�-4FhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ��g�?*;L]n�?*             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJr��<hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�B                          ���?�������?%             N@                         �S�?��Sݭg�?            �C@������������������������       �                     $@������������������������       �                     =@������������������������       ������?             5@�t�bh�h(h+K ��h-��R�(KKKK��hW�CP      =@      ?@      $@      =@      $@                      =@      3@       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�D�thG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?*;L]n�?'             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�o7hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�B                          `;0�?d��0u��?#             N@������������������������       �        	             2@                         �L�?�G��l��?             E@������������������������       �                     6@������������������������       �        
             4@�t�bh�h(h+K ��h-��R�(KKKK��hW�CP      6@      C@              2@      6@      4@      6@                      4@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ"�hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?��S���?*             N@������������������������       �                     <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      <@      @@      <@                      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���"hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?d��0u��?$             N@������������������������       �                    �B@������������������������       ��nkK�?             7@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      C@      6@     �B@              �?      6@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�h�hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��q�q�?)             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      4@      D@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���RhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?�������?&             N@������������������������       �                     =@������������������������       �                     ?@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      =@                      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ5\hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?��S���?)             N@������������������������       �                     :@������������������������       ��IєX�?             A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      <@      @@      :@               @      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�Q&hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�������?'             N@������������������������       �      �?             @@������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ?@      =@      ?@      �?              <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ&N�hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��G�z��?+             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      ;@     �@@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��8hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?�������?*             N@������������������������       �                     =@������������������������       �                     ?@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      =@                      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�b�hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?      �?"             N@������������������������       ��g�y��?             ?@������������������������       �                     =@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      >@      >@      >@      �?              =@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��bhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?��Q��?*             N@������������������������       �                     5@������������������������       �                    �C@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      5@     �C@      5@                     �C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJOy�qhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�G�z��?"             N@������������������������       �                     ;@������������������������       �                    �@@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ;@     �@@      ;@                     �@@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��ghG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?      �?%             N@������������������������       �                     <@������������������������       �      �?             @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      >@      >@      <@               @      >@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJiƋ.hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        p���?�G�z��?             N@������������������������       �`Jj��?             ?@������������������������       �\-��p�?             =@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      ;@     �@@       @      =@      9@      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ*�/shG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?��S���?'             N@������������������������       �                     @@������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      @@      <@      @@                      <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��\hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       �*;L]n�?'             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      :@      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�B                          `;0�?�������?#             N@������������������������       ������H�?
             2@                         ���?X�Cc�?             E@������������������������       �                     ;@������������������������       �                     .@�t�bh�h(h+K ��h-��R�(KKKK��hW�CP      =@      ?@       @      0@      ;@      .@      ;@                      .@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJxS�ohG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?��S���?&             N@������������������������       �                     <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      <@      @@      <@                      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJQ ghG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        ����?��Q��?%             N@������������������������       �                     5@������������������������       �                    �C@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      5@     �C@      5@                     �C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJA��2hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?*;L]n�?&             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ojhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         @>��?d��0u��?*             N@������������������������       �                     6@������������������������       �                     C@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      6@      C@      6@                      C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��jhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�q�q�?#             N@������������������������       � ��WV�?             :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      9@     �A@      9@      �?              A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ9hExhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?��S���?!             N@������������������������       �                     <@������������������������       �                     @@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      <@      @@      <@                      @@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ#9�*hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��q�q�?'             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C     �A@      9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJf/4'hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         ���?      �?(             N@������������������������       �                     >@������������������������       �                     >@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      >@      >@      >@                      >@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJw�+hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                         x��?*;L]n�?*             N@������������������������       �                     :@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@                      A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��+hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�0u��A�?'             N@������������������������       � �q�q�?             8@������������������������       �                     B@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      7@     �B@      7@      �?              B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���5hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��������?)             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      =@      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJRܯ[hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ���S���?"             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      @@      <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ[P!hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?*;L]n�?+             N@������������������������       � 7���B�?             ;@������������������������       �                    �@@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      :@      A@      :@      �?             �@@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��,@hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hK hnKhoh(h+K ��h-��R�(KK��hv�C8������������������������       ��0u��A�?(             N@�t�bh�h(h+K ��h-��R�(KKKK��hW�C      7@     �B@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��PhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        �$I�?�������?)             N@������������������������       �`Jj��?             ?@������������������������       �                     =@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      =@       @              =@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJcʚhG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�������?&             N@������������������������       �                     =@������������������������       �                     ?@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0      =@      ?@      =@                      ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ5&]hG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                        жm�?�q�q�?!             N@������������������������       �                     A@������������������������       � ��WV�?             :@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0     �A@      9@      A@              �?      9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�K6ShG        hNhG?��G�z�h=Kh>Kh?h(h+K ��h-��R�(KK��hW�C              �?�t�bhKh\hFC       ���R�h`KhahdKh(h+K ��h-��R�(KK��hF�C       �t�bK��R�}�(hKhnKhoh(h+K ��h-��R�(KK��hv�C�                           �?�0u��A�?(             N@������������������������       �                    �B@������������������������       �                     7@�t�bh�h(h+K ��h-��R�(KKKK��hW�C0     �B@      7@     �B@                      7@�t�bubhhubehhub.